library verilog;
use verilog.vl_types.all;
entity Extend_Unit_tb is
end Extend_Unit_tb;
