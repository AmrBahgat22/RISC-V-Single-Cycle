library verilog;
use verilog.vl_types.all;
entity Program_Counter_tb is
end Program_Counter_tb;
